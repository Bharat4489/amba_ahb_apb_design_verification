module ahb_arbiter (
    ahb_if.arbiter_mp arbiter_if
);

endmodule